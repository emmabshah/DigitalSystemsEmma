module task210_challenge;
